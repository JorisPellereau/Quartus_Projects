
module nios_leds (
	clk_clk,
	pio_green_leds_0_external_connection_export,
	reset_reset_n);	

	input		clk_clk;
	output	[8:0]	pio_green_leds_0_external_connection_export;
	input		reset_reset_n;
endmodule
