-- altera_vjtag_24ir.vhd

-- Generated using ACDS version 20.1 720

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity altera_vjtag_24ir is
	port (
		tdi                : out std_logic;                                        -- jtag.tdi
		tdo                : in  std_logic                     := '0';             --     .tdo
		ir_in              : out std_logic_vector(23 downto 0);                    --     .ir_in
		ir_out             : in  std_logic_vector(23 downto 0) := (others => '0'); --     .ir_out
		virtual_state_cdr  : out std_logic;                                        --     .virtual_state_cdr
		virtual_state_sdr  : out std_logic;                                        --     .virtual_state_sdr
		virtual_state_e1dr : out std_logic;                                        --     .virtual_state_e1dr
		virtual_state_pdr  : out std_logic;                                        --     .virtual_state_pdr
		virtual_state_e2dr : out std_logic;                                        --     .virtual_state_e2dr
		virtual_state_udr  : out std_logic;                                        --     .virtual_state_udr
		virtual_state_cir  : out std_logic;                                        --     .virtual_state_cir
		virtual_state_uir  : out std_logic;                                        --     .virtual_state_uir
		tck                : out std_logic                                         --  tck.clk
	);
end entity altera_vjtag_24ir;

architecture rtl of altera_vjtag_24ir is
	component sld_virtual_jtag is
		generic (
			sld_auto_instance_index : string  := "YES";
			sld_instance_index      : integer := 0;
			sld_ir_width            : integer := 1
		);
		port (
			tdi                : out std_logic;                                        -- tdi
			tdo                : in  std_logic                     := 'X';             -- tdo
			ir_in              : out std_logic_vector(23 downto 0);                    -- ir_in
			ir_out             : in  std_logic_vector(23 downto 0) := (others => 'X'); -- ir_out
			virtual_state_cdr  : out std_logic;                                        -- virtual_state_cdr
			virtual_state_sdr  : out std_logic;                                        -- virtual_state_sdr
			virtual_state_e1dr : out std_logic;                                        -- virtual_state_e1dr
			virtual_state_pdr  : out std_logic;                                        -- virtual_state_pdr
			virtual_state_e2dr : out std_logic;                                        -- virtual_state_e2dr
			virtual_state_udr  : out std_logic;                                        -- virtual_state_udr
			virtual_state_cir  : out std_logic;                                        -- virtual_state_cir
			virtual_state_uir  : out std_logic;                                        -- virtual_state_uir
			tck                : out std_logic                                         -- clk
		);
	end component sld_virtual_jtag;

begin

	virtual_jtag_0 : component sld_virtual_jtag
		generic map (
			sld_auto_instance_index => "NO",
			sld_instance_index      => 0,
			sld_ir_width            => 24
		)
		port map (
			tdi                => tdi,                -- jtag.tdi
			tdo                => tdo,                --     .tdo
			ir_in              => ir_in,              --     .ir_in
			ir_out             => ir_out,             --     .ir_out
			virtual_state_cdr  => virtual_state_cdr,  --     .virtual_state_cdr
			virtual_state_sdr  => virtual_state_sdr,  --     .virtual_state_sdr
			virtual_state_e1dr => virtual_state_e1dr, --     .virtual_state_e1dr
			virtual_state_pdr  => virtual_state_pdr,  --     .virtual_state_pdr
			virtual_state_e2dr => virtual_state_e2dr, --     .virtual_state_e2dr
			virtual_state_udr  => virtual_state_udr,  --     .virtual_state_udr
			virtual_state_cir  => virtual_state_cir,  --     .virtual_state_cir
			virtual_state_uir  => virtual_state_uir,  --     .virtual_state_uir
			tck                => tck                 --  tck.clk
		);

end architecture rtl; -- of altera_vjtag_24ir
